library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity MaquinaEstado is
Port ( CLK : in STD_LOGIC;
           BTN : in STD_LOGIC_VECTOR (4 downto 0);
           LED : out STD_LOGIC_VECTOR (15 downto 0));
end MaquinaEstado;

architecture Behavioral of MaquinaEstado is

begin


end Behavioral;

